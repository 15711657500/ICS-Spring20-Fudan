module conflict (
    input logic branchD, memtoregE, regwriteE, memtoregM, regwriteM, regwriteW,
    input logic [4:0]rsD, rtD, rsE, rtE, writeregE, writeregM, writeregW,
    output logic stallF, stallD, forwardAD, forwardBD, flushE, forwardAE, forwardBE
);
    
endmodule